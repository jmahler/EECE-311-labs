EECE 311 Example 1

VS 0 1 DC 100V
IS 0 3 DC 5A
R1 1 2 10
R2 2 5 20
R3 3 0 50
R4 3 4 40
E1 4 0 1 0 0.5
F1 0 2 VS 0.5
G1 4 3 1 0 0.1
H1 1 3 VX 2
VX 5 3 DC 0V

.DC VS 0V 100V 5V
.PRINT DC I(R1) I(R2) I(R3) I(R4)
.PRINT DC V(1) V(2) V(3) V(4) V(5)
.PLOT DC V(0,4)
.PROBE
.END
