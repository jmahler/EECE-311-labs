EECE 311 Laboratory Project #2
* run using: ngspice -b lab1.cir
* http://www.ecst.csuchico.edu/~hma/Lab2.311.pdf

VS1 10 0 DC 50V
VSENS 10 1 DC 0V
R1 1 2 6
R2 0 2 8
R3 2 3 2
R4 0 3 4
* current controlled current source
F1 2 3 VSENS 3
I1 0 3 DC 5

* sweep VS1 from 0 volts to 50 volts in 10 volt increments
.DC VS1 0V 50V 10V

.PRINT DC V(2) V(3)
*.PLOT DC V(1) V(2) V(3)
.PRINT DC I(VS1) I(F1) I(R1) I(R2) I(R3) I(R4)

*.PROBE
.END