EECE 311, Lab 4, example 2: pulsed response RLC circuit

* PWL( t0 v0 t1 v1 t2 v2)
V1 1 0 PWL(0 0 1NS 1V 1MS 1V)

R1 1 2 2
L1 2 3 50uH
C1 3 0 10uF

V2 4 0 PWL(0 0 1NS 1V 1MS 1V)
R2 4 5 1
L2 5 6 50uH
C2 6 0 10uF

V3 7 0 PWL(0 0 1NS 1V 1MS 1V)
R3 7 8 8
L3 8 9 50uH
C3 9 0 10uF

* .TRAN step end_time
.TRAN 1uS 500uS
.PLOT TRAN V(3) V(6) V(9)
.PROBE

.END